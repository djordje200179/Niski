localparam INST_LUI				= 7'b0110111,
		   INST_AUIPC		   	= 7'b0010111,
		   INST_JAL			 	= 7'b1101111,
		   INST_JALR			= 7'b1100111,
		   INST_GROUP_BRANCH	= 7'b1100011,
		   INST_GROUP_LOAD		= 7'b0000011,
		   INST_GROUP_STORE		= 7'b0100011,
		   INST_GROUP_ARLOG_IMM	= 7'b0010011,
		   INST_GROUP_ARLOG		= 7'b0110011,
		   INST_GROUP_MISC_MEM	= 7'b0001111,
		   INST_GROUP_SYSTEM	= 7'b1110011;

localparam INST_BRANCH_EQ   = 3'b000,
		   INST_BRANCH_NEQ  = 3'b001,
		   INST_BRANCH_LT   = 3'b100,
		   INST_BRANCH_GE   = 3'b101,
		   INST_BRANCH_LTU  = 3'b110,
		   INST_BRANCH_GEU  = 3'b111;

localparam INST_LOAD_BYTE	   	= 3'b000,
		   INST_LOAD_HALF	   	= 3'b001,
		   INST_LOAD_WORD	   	= 3'b010,
		   INST_LOAD_BYTE_UNS 	= 3'b100,
		   INST_LOAD_HALF_UNS	= 3'b101;

localparam INST_STORE_BYTE	  = 3'b000,
		   INST_STORE_HALF	  = 3'b001,
		   INST_STORE_WORD	  = 3'b010;

localparam INST_ARLOG_ADD	= 3'b000,
		   INST_ARLOG_SL 	= 3'b001,
		   INST_ARLOG_SLT 	= 3'b010,
		   INST_ARLOG_SLTU	= 3'b011,
		   INST_ARLOG_XOR 	= 3'b100,
		   INST_ARLOG_SR 	= 3'b101,
		   INST_ARLOG_OR 	= 3'b110,
		   INST_ARLOG_AND 	= 3'b111;

localparam INST_ADD_MOD_ADD = 7'b0000000,
		   INST_ADD_MOD_SUB = 7'b0100000;

localparam INST_SR_MOD_L = 7'b0000000,
		   INST_SR_MOD_A = 7'b0100000;

// TODO: Add for FENCE, FENCE.TSO, PAUSE

localparam INST_SYSTEM_ECALL 	= 12'b000000000000,
		   INST_SYSTEM_EBREAK 	= 12'b000000000001;