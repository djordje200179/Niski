localparam PS2_KEYBOARD_BRK_CODE = 8'hF0,
		   PS2_KEYBOARD_EXT_CODE = 8'hE0,
		   
		   PS2_KEYBOARD_NUMPAD_0 = 8'h70,
		   PS2_KEYBOARD_NUMPAD_1 = 8'h69,
		   PS2_KEYBOARD_NUMPAD_2 = 8'h72,
		   PS2_KEYBOARD_NUMPAD_3 = 8'h7A,
		   PS2_KEYBOARD_NUMPAD_4 = 8'h6B,
		   PS2_KEYBOARD_NUMPAD_5 = 8'h73,
		   PS2_KEYBOARD_NUMPAD_6 = 8'h74,
		   PS2_KEYBOARD_NUMPAD_7 = 8'h6C,
		   PS2_KEYBOARD_NUMPAD_8 = 8'h75,
		   PS2_KEYBOARD_NUMPAD_9 = 8'h7D,
		   
		   PS2_KEYBOARD_NUMPAD_E_DIV= 8'h4A,
		   PS2_KEYBOARD_NUMPAD_MUL	= 8'h7C,
		   PS2_KEYBOARD_NUMPAD_MIN 	= 8'h7B,
		   PS2_KEYBOARD_NUMPAD_PLUS = 8'h79,
		   
		   PS2_KEYBOARD_0 = 8'h45,
		   PS2_KEYBOARD_1 = 8'h16,
		   PS2_KEYBOARD_2 = 8'h1E,
		   PS2_KEYBOARD_3 = 8'h26,
		   PS2_KEYBOARD_4 = 8'h25,
		   PS2_KEYBOARD_5 = 8'h2E,
		   PS2_KEYBOARD_6 = 8'h36,
		   PS2_KEYBOARD_7 = 8'h3D,
		   PS2_KEYBOARD_8 = 8'h3E,
		   PS2_KEYBOARD_9 = 8'h46,
		   
		   PS2_KEYBOARD_ENTER = 8'h5A,
		   PS2_KEYBOARD_SPACE = 8'h29,
		   
		   PS2_KEYBOARD_E_LEFT	= 8'h6B,
		   PS2_KEYBOARD_E_UP	= 8'h75,
		   PS2_KEYBOARD_E_RIGHT	= 8'h74,
		   PS2_KEYBOARD_E_DOWN	= 8'h72;

