`ifndef I2C_STATES
`define I2C_STATES

localparam STATE_IDLE = 3'd0;

`endif