localparam STATE_IDLE	= 2'd0,
		   STATE_CPU	= 2'd1,
		   STATE_DMA	= 2'd2;